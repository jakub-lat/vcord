module models

pub struct User {
	pub:
	username string
	discriminator string
}