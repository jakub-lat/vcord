module config

import vcord.utils

pub struct Config {
pub:
	token	string
	log_level utils.LogLevel
}