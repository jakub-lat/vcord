module models

struct User {
	id					string
}