module vcord

// TODO