module main

import vcord

fn main() {
	_ := vcord.create_client()
}
