module models

const (
	create_instant_invite = 1 << 0
	kick_members = 1 << 1
	ban_members = 1 << 2
	administrator = 1 << 3
	manage_channels = 1 << 4
	manage_guild = 1 << 5
	add_reactions = 1 << 6
	view_audit_log = 1 << 7
	priority_speaker = 1 << 8
	stream = 1 << 9
	view_channel = 1 << 10
	send_messages = 1 << 11
	send_tts_messages = 1 << 12
	manage_messages = 1 << 13
	embed_links = 1 << 14
	attach_files = 1 << 15
	read_message_history = 1 << 16
	mention_everyone = 1 << 17
	use_external_emojis = 1 << 18
	view_guild_insights = 1 << 19
	connect = 1 << 20
	speak = 1 << 21
	mute_members = 1 << 22
	deafen_members = 1 << 23
	move_members = 1 << 24
	use_voice_activity = 1 << 25
	change_nickname = 1 << 26
	manage_nicknames = 1 << 27
	manage_roles = 1 << 28
	manage_webhooks = 1 << 29
	manage_emojis = 1 << 30
)

type Perms int

pub fn parse_perms(i int) Perms {
	return Perms(i)
}